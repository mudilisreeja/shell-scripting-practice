id,name,age
01,paul,20
02,alex,30
03,raju,4
	
